
// this is where things get wild...
module neuron #(parameter bias_file="", weight_file="", num_of_weights=764);

// loading the data from memory. This will be a signifigent challenge. 
	// might include some nested terenary operators...

// memory
	// note, r_address is incrimented up by one each "loop".



endmodule
