

module adder_tb;
reg [31:0] x;
reg [31:0] y;
reg c_in;
wire c_out;
wire [31:0] sum;

adder a (.x(x), .y(y), .c_in(c_in), .c_out(c_out), .sum(sum));

initial begin

x = 32'b0000000000000000_0000000000000000;
y = 32'b0000000000000000_0000000000000001;
c_in = 0;
#20
x = 32'b0000000000000000_0000000000000001;
y = 32'b0000000000000000_0000000000000001;
c_in = 1;
#20
x = 32'b1000000000000000_0000000000000000;
y = 32'b1000000000000000_0000000000000001;
c_in = 0;
#20
x = 32'b0000000000000000_0000111110000001;
y = 32'b0000000000000000_0000000011110001;
c_in = 0;

end 

endmodule	
